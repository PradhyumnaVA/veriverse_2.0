module first_prog();

initial begin
	$display("hello world");
end

endmodule
